library ieee;
use ieee.std_logic_1164.all;

entity counter is
port (
    clk_i       : in  std_logic;
    rst_i       : in  std_logic;
    -- TODO : Add in and out ports
);
end counter;

