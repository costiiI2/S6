library ieee;
use ieee.std_logic_1164.all;

package counterg_pkg is

      type counter_in_type is record
      	-- TODO : Complete
      end record;

      type counter_out_type is record
      	-- TODO : Complete
      end record;

end package;
